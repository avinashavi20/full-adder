/********************************************************************************************

Copyright 2018-2019 - Maven Silicon Softech Pvt Ltd. All Rights Reserved.

This source code is an unpublished work belongs to Maven Silicon Softech Pvt Ltd.
It is considered a trade secret and is not to be divulged or used by parties who 
have not received written authorization from Maven Silicon Softech Pvt Ltd.

Maven Silicon Softech Pvt Ltd
Bangalore - 560076

Webpage: www.maven-silicon.com

Filename:	full_adder.v   

Description:	One bit Full adder design 

Date:		01/05/2018

Author:		Maven Silicon

Email:		online@maven-silicon.com
			 

Version:	1.0

*********************************************************************************************/

module full_adder(a,
                  b,
                  c,
                  sum,
                  carry);

  // Step 1. Write down the directions for the ports	     

input a,b,c;
output sum, carry;

assign sum = a ^ b ^ c;
assign carry = a & b | b & c | c & a;
  // Step 2. Declare the internal wires    


  // Step 3. Instantiate two Half-Adders


  // Step 4. Instantiate the OR gate


endmodule

